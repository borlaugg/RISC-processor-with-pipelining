library ieee;
use ieee.std_logic_1164.all;
package Decoderpkg is
	component decoder is
		port(instruction:in std_logic_vector(15 downto 0);
			  cz:in std_logic_vector(1 downto 0);
			  bp,clock:in std_logic;
			  yz: out std_logic_vector(1 downto 0);
			  imm6: out std_logic_vector(5 downto 0);
			  rf_rs, rf_ws: out std_logic_vector(7 downto 0);
			  imm9: out std_logic_vector(8 downto 0);
			  c_we, c_re, z_we, z_re, d_re0, d_we0,d_re1, d_we1,d_re2, d_we2,d_re3, 
			  d_we3,d_re4, d_we4,d_re5, d_we5,d_re6, d_we6,d_we7,d_re7: out std_logic;
			  opcode: out std_logic_vector(3 downto 0));
	end component decoder;
end package Decoderpkg;

library ieee;
use ieee.std_logic_1164.all;
library work;
use work.DecodeRegpkg.all;

entity decoder is
	port(instruction:in std_logic_vector(15 downto 0);
		  cz:in std_logic_vector(1 downto 0);
		  bp,clock:in std_logic;
		  yz: out std_logic_vector(1 downto 0);
		  imm6: out std_logic_vector(5 downto 0);
		  rf_rs, rf_ws: out std_logic_vector(7 downto 0);
		  imm9: out std_logic_vector(8 downto 0);
		  c_we, c_re, z_we, z_re, d_re0, d_we0,d_re1, d_we1,d_re2, d_we2,d_re3, 
		  d_we3,d_re4, d_we4,d_re5, d_we5,d_re6, d_we6,d_we7,d_re7: out std_logic;
		  opcode: out std_logic_vector(3 downto 0));
end decoder;

architecture beh of decoder is
signal op : std_logic_vector(3 downto 0);
signal rfa,rfb,rfc: std_logic_vector(7 downto 0);
signal xy : std_logic_vector(1 downto 0);
signal ra, rb, rc : std_logic_vector(2 downto 0);
begin
op <= instruction (15 downto 12);
xy <=	instruction (1 downto 0);
ra <=	instruction (11 downto 9);
rb <=	instruction (8 downto 6);
rc <=	instruction (5 downto 3); 
dec1: DecodeReg port map(ra => ra, rf => rfa);
dec2: DecodeReg port map(ra => rb, rf => rfb);
dec3: DecodeReg port map(ra => rc, rf => rfc);
decode:process(clock)
	begin	
		if (clock' event and clock= '1' and bp ='0') then
			case op is
				when "0000"=> -- ADDI
					opcode <= op;
					yz <= "00";
					imm6 <= instruction(5 downto 0);
					imm9 <="000000000";
					c_we <= '1';
					z_we <= '1';
					c_re <= '0';
					z_re <= '0';
					d_re0 <= '0';
					d_we0 <= '0';
					d_re1 <= '0';
					d_we1 <= '0';
					d_re2 <= '0';
					d_we2 <= '0';
					d_re3 <= '0'; 
					d_we3 <= '0';
					d_re4 <= '0';
					d_we4 <= '0';
					d_re5 <= '0'; 
					d_we5 <= '0';
					d_re6 <= '0'; 
					d_we6 <= '0';
					d_re7 <= '0'; 
					d_we7 <= '0';	
					rf_rs <= rfb;
					rf_ws <= rfa;
				when "0001"=> -- ADD
					opcode <= op;
					yz <= xy;
					imm6 <= "000000";
					imm9 <="000000000";
					c_we <= '1';
					z_we <= '1';
					c_re <= '0';
					z_re <= '0';
					d_re0 <= '0';
					d_we0 <= '0';
					d_re1 <= '0';
					d_we1 <= '0';
					d_re2 <= '0';
					d_we2 <= '0';
					d_re3 <= '0'; 
					d_we3 <= '0';
					d_re4 <= '0';
					d_we4 <= '0';
					d_re5 <= '0'; 
					d_we5 <= '0';
					d_re6 <= '0'; 
					d_we6 <= '0'; 
					d_re7 <= '0'; 
					d_we7 <= '0';
					if( xy = "00") then
						rf_rs(0) <= rfb(0) or rfc(0);
						rf_rs(1) <= rfb(1) or rfc(1);
						rf_rs(2) <= rfb(2) or rfc(2);
						rf_rs(3) <= rfb(3) or rfc(3);
						rf_rs(4) <= rfb(4) or rfc(4);
						rf_rs(5) <= rfb(5) or rfc(5);
						rf_rs(6) <= rfb(6) or rfc(6);
						rf_rs(7) <= rfb(7) or rfc(7);
						rf_ws <= rfa;
					elsif( xy = "10") then 
						if( cz(0) = '1') then
							rf_rs(0) <= rfb(0) or rfc(0);
							rf_rs(1) <= rfb(1) or rfc(1);
							rf_rs(2) <= rfb(2) or rfc(2);
							rf_rs(3) <= rfb(3) or rfc(3);
							rf_rs(4) <= rfb(4) or rfc(4);
							rf_rs(5) <= rfb(5) or rfc(5);
							rf_rs(6) <= rfb(6) or rfc(6);
							rf_rs(7) <= rfb(7) or rfc(7);
							rf_ws <= rfa;
						elsif ( cz(0) ='0') then
							rf_rs <= "00000000";
							rf_ws <= "00000000";
						end if;
					elsif( xy = "01") then
						if( cz(1) = '1') then
							rf_rs(0) <= rfb(0) or rfc(0);
							rf_rs(1) <= rfb(1) or rfc(1);
							rf_rs(2) <= rfb(2) or rfc(2);
							rf_rs(3) <= rfb(3) or rfc(3);
							rf_rs(4) <= rfb(4) or rfc(4);
							rf_rs(5) <= rfb(5) or rfc(5);
							rf_rs(6) <= rfb(6) or rfc(6);
							rf_rs(7) <= rfb(7) or rfc(7);
							rf_ws <= rfa;
						elsif ( cz(1) ='0') then
							rf_rs <= "00000000";
							rf_ws <= "00000000";
						end if;
					elsif (xy = "11") then
						rf_rs(0) <= rfb(0) or rfc(0);
						rf_rs(1) <= rfb(1) or rfc(1);
						rf_rs(2) <= rfb(2) or rfc(2);
						rf_rs(3) <= rfb(3) or rfc(3);
						rf_rs(4) <= rfb(4) or rfc(4);
						rf_rs(5) <= rfb(5) or rfc(5);
						rf_rs(6) <= rfb(6) or rfc(6);
						rf_rs(7) <= rfb(7) or rfc(7);
						rf_ws <= rfa;
					end if;
				when "0010"=> -- 	NAND
					opcode <= op;
					yz <= xy;
					imm6 <= "000000";
					imm9 <="000000000";
					c_we <= '0';
					z_we <= '1';
					c_re <= '0';
					z_re <= '0';
					d_re0 <= '0';
					d_we0 <= '0';
					d_re1 <= '0';
					d_we1 <= '0';
					d_re2 <= '0';
					d_we2 <= '0';
					d_re3 <= '0'; 
					d_we3 <= '0';
					d_re4 <= '0';
					d_we4 <= '0';
					d_re5 <= '0'; 
					d_we5 <= '0';
					d_re6 <= '0'; 
					d_we6 <= '0';
					d_re7 <= '0'; 
					d_we7 <= '0';
						if( xy = "00") then
							rf_rs(0) <= rfb(0) or rfc(0);
							rf_rs(1) <= rfb(1) or rfc(1);
							rf_rs(2) <= rfb(2) or rfc(2);
							rf_rs(3) <= rfb(3) or rfc(3);
							rf_rs(4) <= rfb(4) or rfc(4);
							rf_rs(5) <= rfb(5) or rfc(5);
							rf_rs(6) <= rfb(6) or rfc(6);
							rf_rs(7) <= rfb(7) or rfc(7);
							rf_ws <= rfa;
						elsif (xy = "01") then
							if( cz(1) = '1') then
								rf_rs(0) <= rfb(0) or rfc(0);
								rf_rs(1) <= rfb(1) or rfc(1);
								rf_rs(2) <= rfb(2) or rfc(2);
								rf_rs(3) <= rfb(3) or rfc(3);
								rf_rs(4) <= rfb(4) or rfc(4);
								rf_rs(5) <= rfb(5) or rfc(5);
								rf_rs(6) <= rfb(6) or rfc(6);
								rf_rs(7) <= rfb(7) or rfc(7);
								rf_ws <= rfa;
							elsif ( cz(1) ='0') then
								rf_rs <= "00000000";
								rf_ws <= "00000000";
							end if;
						elsif( xy = "10") then
							if( cz(0) = '1') then
								rf_rs(0) <= rfb(0) or rfc(0);
								rf_rs(1) <= rfb(1) or rfc(1);
								rf_rs(2) <= rfb(2) or rfc(2);
								rf_rs(3) <= rfb(3) or rfc(3);
								rf_rs(4) <= rfb(4) or rfc(4);
								rf_rs(5) <= rfb(5) or rfc(5);
								rf_rs(6) <= rfb(6) or rfc(6);
								rf_rs(7) <= rfb(7) or rfc(7);
								rf_ws <= rfa;
							elsif ( cz(0) ='0') then
								rf_rs <= "00000000";
								rf_ws <= "00000000";
							end if;
						else
							rf_rs <= "00000000";
							rf_ws <= "00000000";
					end if;
				when "0101"=> -- SW
					opcode <= op;
					yz <= "00";
					imm6 <= instruction(5 downto 0);
					imm9 <="000000000";
					c_we <= '0';
					z_we <= '0';
					c_re <= '0';
					z_re <= '0';
					d_re0 <= '0';
					d_we0 <= rfa(0);
					d_re1 <= '0';
					d_we1 <= rfa(1);
					d_re2 <= '0';
					d_we2 <= rfa(2);
					d_re3 <= '0'; 
					d_we3 <= rfa(3);
					d_re4 <= '0';
					d_we4 <= rfa(4);
					d_re5 <= '0'; 
					d_we5 <= rfa(5);
					d_re6 <= '0'; 
					d_we6 <= rfa(6);
					d_re7 <= '0'; 
					d_we7 <= rfa(7);
					rf_rs(0) <= rfb(0) or rfa(0);
					rf_rs(1) <= rfb(1) or rfa(1);
					rf_rs(2) <= rfb(2) or rfa(2);
					rf_rs(3) <= rfb(3) or rfa(3);
					rf_rs(4) <= rfb(4) or rfa(4);
					rf_rs(5) <= rfb(5) or rfa(5);
					rf_rs(6) <= rfb(6) or rfa(6);
					rf_rs(7) <= rfb(7) or rfa(7);
					rf_ws <= "00000000";
				when "0111"=> -- LW
					opcode <= op;
					yz <= "00";
					imm6 <= instruction(5 downto 0);
					imm9 <="000000000";
					c_we <= '0';
					z_we <= '0';
					c_re <= '0';
					z_re <= '0';
					d_we0 <= '0';
					d_re0 <= rfa(0);
					d_we1 <= '0';
					d_re1 <= rfa(1);
					d_we2 <= '0';
					d_re2 <= rfa(2);
					d_we3 <= '0'; 
					d_re3 <= rfa(3);
					d_we4 <= '0';
					d_re4 <= rfa(4);
					d_we5 <= '0'; 
					d_re5 <= rfa(5);
					d_we6 <= '0'; 
					d_re6 <= rfa(6);
					d_we7 <= '0'; 
					d_re7 <= rfa(7);
					rf_rs <= rfb;
					rf_ws <= rfa;
				when "1000"=> -- BEQ
					opcode <= op;
					yz <= "00";
					imm6 <= instruction(5 downto 0);
					imm9 <="000000000";
					c_we <= '0';
					z_we <= '0';
					c_re <= '0';
					z_re <= '0';
					d_re0 <= '0';
					d_we0 <= '0';
					d_re1 <= '0';
					d_we1 <= '0';
					d_re2 <= '0';
					d_we2 <= '0';
					d_re3 <= '0'; 
					d_we3 <= '0';
					d_re4 <= '0';
					d_we4 <= '0';
					d_re5 <= '0'; 
					d_we5 <= '0';
					d_re6 <= '0'; 
					d_we6 <= '0';
					d_re7 <= '0'; 
					d_we7 <= '0';
					rf_rs(0) <= rfb(0) or rfa(0);
					rf_rs(1) <= rfb(1) or rfa(1);
					rf_rs(2) <= rfb(2) or rfa(2);
					rf_rs(3) <= rfb(3) or rfa(3);
					rf_rs(4) <= rfb(4) or rfa(4);
					rf_rs(5) <= rfb(5) or rfa(5);
					rf_rs(6) <= rfb(6) or rfa(6);
					rf_rs(7) <= rfb(7) or rfa(7);
					rf_ws <= "00000000";
				when "1001"=> -- JAL
					opcode <= op;
					yz <= "00";
					imm6 <= "000000";
					imm9 <=instruction(8 downto 0);
					c_we <= '0';
					z_we <= '0';
					c_re <= '0';
					z_re <= '0';
					d_re0 <= '0';
					d_we0 <= '0';
					d_re1 <= '0';
					d_we1 <= '0';
					d_re2 <= '0';
					d_we2 <= '0';
					d_re3 <= '0'; 
					d_we3 <= '0';
					d_re4 <= '0';
					d_we4 <= '0';
					d_re5 <= '0'; 
					d_we5 <= '0';
					d_re6 <= '0'; 
					d_we6 <= '0';
					d_re7 <= '0'; 
					d_we7 <= '0';
					rf_rs <= "00000000";
					rf_ws <= rfa;
				when "1010"=> -- JLR
					opcode <= op;
					yz <= "00";
					imm6 <= "000000";
					imm9 <="000000000";
					c_we <= '0';
					z_we <= '0';
					c_re <= '0';
					z_re <= '0';
					d_re0 <= '0';
					d_we0 <= '0';
					d_re1 <= '0';
					d_we1 <= '0';
					d_re2 <= '0';
					d_we2 <= '0';
					d_re3 <= '0'; 
					d_we3 <= '0';
					d_re4 <= '0';
					d_we4 <= '0';
					d_re5 <= '0'; 
					d_we5 <= '0';
					d_re6 <= '0'; 
					d_we6 <= '0';
					d_re7 <= '0'; 
					d_we7 <= '0';
					rf_rs <= rfb;
					rf_ws <= rfa;
				when "1011"=> -- JRI
					opcode <= op;
					yz <= "00";
					imm6 <= "000000";
					imm9 <=instruction(8 downto 0);
					c_we <= '0';
					z_we <= '0';
					c_re <= '0';
					z_re <= '0';
					d_re0 <= '0';
					d_we0 <= '0';
					d_re1 <= '0';
					d_we1 <= '0';
					d_re2 <= '0';
					d_we2 <= '0';
					d_re3 <= '0'; 
					d_we3 <= '0';
					d_re4 <= '0';
					d_we4 <= '0';
					d_re5 <= '0'; 
					d_we5 <= '0';
					d_re6 <= '0'; 
					d_we6 <= '0';
					d_re7 <= '0'; 
					d_we7 <= '0';
					rf_rs <= rfa;
					rf_ws <= "00000000";
				when "1101"=> -- SM
					opcode <= op;
					yz <= "00";
					imm6 <= "000000";
					imm9 <="000000000";
					c_we <= '0';
					z_we <= '0';
					c_re <= '0';
					z_re <= '0';
					d_re0 <= instruction(0);
					d_we0 <= '0';
					d_re1 <= instruction(1);
					d_we1 <= '0';
					d_re2 <= instruction(2);
					d_we2 <= '0';
					d_re3 <= instruction(3); 
					d_we3 <= '0';
					d_re4 <= instruction(4);
					d_we4 <= '0';
					d_re5 <= instruction(5); 
					d_we5 <= '0';
					d_re6 <= instruction(6); 
					d_we6 <= '0'; 
					d_re7 <= instruction(7); 
					d_we7 <= '0';
					rf_rs <= rfa;
					rf_ws <= instruction(7 downto 0);
				when "1111"=> --LHI
					opcode <= op;
					yz <= "00";
					imm6 <= "000000";
					imm9 <=instruction(8 downto 0);
					c_we <= '0';
					z_we <= '0';
					c_re <= '0';
					z_re <= '0';
					d_re0 <= '0';
					d_we0 <= '0';
					d_re1 <= '0';
					d_we1 <= '0';
					d_re2 <= '0';
					d_we2 <= '0';
					d_re3 <= '0'; 
					d_we3 <= '0';
					d_re4 <= '0';
					d_we4 <= '0';
					d_re5 <= '0'; 
					d_we5 <= '0';
					d_re6 <= '0'; 
					d_we6 <= '0';
					d_re7 <= '0'; 
					d_we7 <= '0';	
					rf_rs <= "00000000";
					rf_ws <= rfa;
				when others =>
					opcode <= "0000";
					yz <= "00";
					imm6 <= "000000";
					imm9 <="000000000";
					c_we <= '0';
					z_we <= '0';
					c_re <= '0';
					z_re <= '0';
					d_re0 <= '0';
					d_we0 <= '0';
					d_re1 <= '0';
					d_we1 <= '0';
					d_re2 <= '0';
					d_we2 <= '0';
					d_re3 <= '0'; 
					d_we3 <= '0';
					d_re4 <= '0';
					d_we4 <= '0';
					d_re5 <= '0'; 
					d_we5 <= '0';
					d_re6 <= '0'; 
					d_we6 <= '0';
					d_re7 <= '0'; 
					d_we7 <= '0';	
					rf_rs <= "00000000";
					rf_ws <= "00000000";
			end case;
		end if;
	end process;

end beh;